module porta_xor (
    input a,
    input b,
    output y
);

    
    xor U1 (y, a, b); 

endmodule