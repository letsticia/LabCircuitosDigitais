module porta_or (
    input a,
    input b,
    output y
);

    or U1 (y, a, b);

endmodule