module porta_not (
    input a,
    output y
);

    not U1 (y, a);

endmodule